`define DWIDTH 8
//module missing reset signal, reset is floating
module seq_mac(a, b, out, reset, clk);
	input [`DWIDTH-1:0] a;
	input [`DWIDTH-1:0] b;
	input reset;
	input clk;
	output [`DWIDTH-1:0] out;
	
	reg [2*`DWIDTH-1:0] out_temp;
	wire [`DWIDTH-1:0] mul_out;
	wire [2*`DWIDTH-1:0] add_out;
	
	reg [`DWIDTH-1:0] a_flopped;
	reg [`DWIDTH-1:0] b_flopped;
	
	wire [2*`DWIDTH-1:0] mul_out_temp;
	reg [2*`DWIDTH-1:0] mul_out_temp_reg;//input is signed or unsigned?
	
	always @(posedge clk) begin//wait one clock cycle 
		if (reset)begin
			a_flopped <= 0;
			b_flopped <= 0;
		end
		else begin
			a_flopped <= a;
			b_flopped <= b;
		end
	end
	
	//assign mul_out = a * b;
	qmult mult_u1(.i_multiplicand(a_flopped), .i_multiplier(b_flopped), .o_result(mul_out_temp));
	
	always @(posedge clk) begin
		if(reset)
			mul_out_temp_reg <= 0;
		else begin
			mul_out_temp_reg <= mul_out_temp;
		end
	end
	
	//we just truncate the higher bits of the product
	//assign add_out = mul_out + out;
	qadd add_u1(.a(out_temp), .b(mul_out_temp_reg), .c(add_out));
	
	always @(posedge clk) begin
		if(reset)
			out_temp <= 0;
		else begin
			out_temp <= add_out;
		end
	end
	
	//down cast the result
	assign out = 
		(out_temp[2*`DWIDTH-1] == 0) ?  //positive number
			(
			   (|(out_temp[2*`DWIDTH-2 : `DWIDTH-1])) ?  //is any bit from 14:7 is 1, that means overlfow
				 {out_temp[2*`DWIDTH-1] , {(`DWIDTH-1){1'b1}}} : //sign bit and then all 1s
				 {out_temp[2*`DWIDTH-1] , out_temp[`DWIDTH-2:0]} 
			)
			: //negative number
			(
			   (|(out_temp[2*`DWIDTH-2 : `DWIDTH-1])) ?  //is any bit from 14:7 is 0, that means overlfow
				 {out_temp[2*`DWIDTH-1] , out_temp[`DWIDTH-2:0]} :// seems wrong?
				 {out_temp[2*`DWIDTH-1] , {(`DWIDTH-1){1'b0}}} //sign bit and then all 0s
			);
	
	endmodule